module NOT_gate (
    input wire a,
    input wire b
);
    
assign b = !a;

endmodule
